library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity rom is
   port( clk      : in std_logic;
         endereco : in unsigned(6 downto 0);
         dado     : out unsigned(15 downto 0) 
   );
end entity;
architecture a_rom of rom is
   type mem is array (0 to 127) of unsigned(15 downto 0);
   constant conteudo_rom : mem := (

      -- caso endereco => conteudo
      0 => B"0100_011_000000000", --LD R3, 0
      1 => B"0100_100_000000000", --LD R4, 0
      2 => B"0001_011_000000000", --MOV A,R3
      3 => B"0111_100_000000000", --ADD A,R4
      4 => B"0010_100_000000000", --MOV R4,A
      5 => B"0011_000_000000001", --LD A,1
      6 => B"0111_011_000000000", --ADD A,R3
      7 => B"0010_011_000000000", --MOV R3,A
      8 => B"0011_000_000011110", --LD A,30
      9 => B"1000_011_000000000", --sub R3,A
      10 => B"0110_001_011111000", --JPB 1, -8
      11 => B"0001_100_000000000", --MOV A,R4
      12 => B"0010_101_000000000", --MOV R5,A
      13 => B"0000_000_000000000", --NOP
   

    --LAB 7
    --0 => B"011111111_001_1111", --LW R1, 0x00FF
    --1 => B"111111111_010_1111", --LD R2, 0x01FF
    --2 => B"010101111_011_1111", --LD R3, 0x00AF
    --3 => B"000011110_100_1111", --LD R4, 0x001E
    --4 => B"101011000_101_1111", --LD R5, 0x0158
    --5 => B"000000000_000_0000", --NOP
    --6 => B"000100001_110_1111", --LD R6, 0x0021
    --7 => B"000000000_000_0000", --NOP
    --8 => B"000101001_111_1111", --LD R7, 0x0029
    --9 => B"000000111_001_0111", --SW R1, R7
    --10 => B"000101010_111_1111", --LD R7, 0x002A
    --11 => B"000000111_010_0111", --SW R2, R7
    --12 => B"000101100_111_1111", --LD R7, 0x002C
    --13 => B"000000111_011_0111", --SW R3, R7
    --14 => B"000101111_111_1111", --LD R7, 0x002F
    --15 => B"000000111_100_0111", --SW R4, R7
    --16 => B"000110101_111_1111", --LD R7, 0x0035
    --17 => B"000000111_101_0111", --SW R5, R7
    --18 => B"000000000_000_0000", --NOP
    --19 => B"000000000_001_1111", --LD R1, 0x0000
    --20 => B"000000000_000_0000", --NOP
    --21 => B"000000001_000_1110", --LD A, 0x0001
    --22 => B"000000000_110_0100", --ADD A, R6
    --23 => B"000000000_110_0010", --MOV R6, A
    --24 => B"000000110_001_1000", --LW R1, R6
    --25 => B"000000000_000_1101", --CLR Z
    --26 => B"000110101_000_1110", --LD A, 0x0035
    --27 => B"000000000_110_0101", --SUB A, R6
    --28 => B"111111001_111_1100", --BNE 0xF9
    --29 => B"000000000_000_0000", --NOP
    --30 => B"000000000_001_0011", --MOV A, R1
    --31 => B"000000000_011_0100", --ADD A, R3
    --32 => B"000000000_100_0010", --MOV R4, A
         
      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture;

